
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package image_pack is
    subtype data_type is std_logic_vector(3 downto 0);

end image_pack;
